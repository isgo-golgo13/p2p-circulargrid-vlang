module node_payload

struct Payload {
    node_id int
    message string
}
