module db

struct Payload {
    id          int
    node_id     int
    payload     string
    received_at string
}
